    Mac OS X            	   2  �     �                                    ATTR;���  �   �  	                  �     com.apple.TextEncoding      �  �  %com.apple.metadata:kMDItemWhereFroms utf-8;134217984bplist00�_�https://udeaeduco.sharepoint.com/sites/LaboratorioCircuitosDigitalesI/_layouts/15/download.aspx?UniqueId=2ef52355-2af9-46f4-9982-36b08b5ae7a7&Translate=false&tempauth=eyJ0eXAiOiJKV1QiLCJhbGciOiJub25lIn0.eyJhdWQiOiIwMDAwMDAwMy0wMDAwLTBmZjEtY2UwMC0wMDAwMDAwMDAwMDAvdWRlYWVkdWNvLnNoYXJlcG9pbnQuY29tQDk5ZTFlNzIxLTcxODQtNDk4ZS04YWZmLWIyYWQ0ZTUzYzFjMiIsImlzcyI6IjAwMDAwMDAzLTAwMDAtMGZmMS1jZTAwLTAwMDAwMDAwMDAwMCIsIm5iZiI6IjE2NTg4Njg0NDgiLCJleHAiOiIxNjU4ODY4NzQ4IiwiZW5kcG9pbnR1cmwiOiJCa09TOFRZNGJXQlgyb2JTRWYra0ZNbjB2K3IyYkYwcXViN0N3cmRGdkpvPSIsImVuZHBvaW50dXJsTGVuZ3RoIjoiMTU3IiwiaXNsb29wYmFjayI6IlRydWUiLCJjaWQiOiJNRGxsTnpVMFlUQXRNVEF5T0Mxa01EQXdMVFEzT0dNdE4yRXpaVGc1T1dVek1XRmsiLCJ2ZXIiOiJoYXNoZWRwcm9vZnRva2VuIiwic2l0ZWlkIjoiTlRJNU1qUXpZemN0WkdWa055MDBPV1ppTFdGaE5Ua3ROakZtTkdRMFpEWTJaV1UzIiwiYXBwX2Rpc3BsYXluYW1lIjoiTWljcm9zb2Z0IFRlYW1zIFdlYiBDbGllbnQiLCJnaXZlbl9uYW1lIjoiSk9TRSIsInNpZ25pbl9zdGF0ZSI6IltcImttc2lcIl0iLCJhcHBpZCI6IjVlM2NlNmMwLTJiMWYtNDI4NS04ZDRiLTc1ZWU3ODc4NzM0NiIsInRpZCI6Ijk5ZTFlNzIxLTcxODQtNDk4ZS04YWZmLWIyYWQ0ZTUzYzFjMiIsInVwbiI6Impvc2UuYWVkb0B1ZGVhLmVkdS5jbyIsInB1aWQiOiIxMDAzM0ZGRkFGNDc4QTU3IiwiY2FjaGVrZXkiOiIwaC5mfG1lbWJlcnNoaXB8MTAwMzNmZmZhZjQ3OGE1N0BsaXZlLmNvbSIsInNjcCI6Im15ZmlsZXMud3JpdGUgYWxsc2l0ZXMuZnVsbGNvbnRyb2wgYWxsc2l0ZXMubWFuYWdlIGFsbHByb2ZpbGVzLndyaXRlIiwidHQiOiIyIiwidXNlUGVyc2lzdGVudENvb2tpZSI6bnVsbCwiaXBhZGRyIjoiMjAwLjI0LjE2LjIzMCJ9.dmt6Y0JaSmMzVGt6SVJFY2Z3d1UrYnd3NjI0VWQ0Z1g4NmlKNlFPcVFsST0&ApiVersion=2.0_https://teams.microsoft.com/  �                           �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          This resource fork intentionally left blank                                                                                                                                                                                                                            ��